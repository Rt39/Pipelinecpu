
module RegDst_mux(
    input [1:0] RegDst,
    input [4:0] RtAddr,
    input [4:0] RdAddr,
    output reg [4:0] RegWriteAddr
);
	always@(RegDst or RtAddr or RdAddr)begin
		case(RegDst)
			2'b00: RegWriteAddr = RtAddr;
			2'b01: RegWriteAddr = RdAddr;
            2'b10: RegWriteAddr = 5'b11111;//$ra 
		endcase
	end
endmodule

module mux2_32(
	input control,
	input [31:0] data0,
	input [31:0] data1,
	output [31:0] out
);
    assign out=control?data1:data0;
endmodule

module DatatoReg_mux(
	input [1:0] DatatoReg,
	input [31:0] ALU_data,
	input [31:0] Mem_data,
	input [31:0] oldPc,
	output reg [31:0] DatatoReg_out
);
	
	always@(ALU_data or Mem_data or DatatoReg)
    begin
		case(DatatoReg)
			2'b00: DatatoReg_out = ALU_data;
			2'b01: DatatoReg_out = Mem_data;
            2'b10: DatatoReg_out = oldPc + 32'd4;
		endcase
	end
endmodule

module Forward_3mux(
    input [31:0] data00,
    input [31:0] data01,
    input [31:0] data10,
    input [1:0] control,
    output [31:0] out
);
    reg [31:0] temp;

    always @(*)
    begin
        case (control)
            2'b00: temp = data00;
            2'b01: temp = data01;
            2'b10: temp = data10;
        endcase
    end
    assign out=temp;
endmodule